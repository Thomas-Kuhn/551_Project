/******************************************************
* Fall 2015 ECE551 Project
* 5-channel Stereo Equalizer
******************************************************/
module Equalizer(clk,RST_n,LED,A2D_SS_n,A2D_MOSI,A2D_SCLK,A2D_MISO,MCLK,SCL,LRCLK,SDout,SDin,AMP_ON,RSTn);

input clk,RST_n;		// 50MHz clock and asynch active low reset from push button
output reg [7:0] LED;		// Active high outputs that drive LEDs
output reg A2D_SS_n;		// Active low slave select to ADC
output reg A2D_MOSI;		// Master Out Slave in to ADC
output reg A2D_SCLK;		// SCLK on SPI interface to ADC
input A2D_MISO;			// Master In Slave Out from ADC
output reg MCLK;			// 12.5MHz clock to CODEC
output reg SCL;				// serial shift clock clock to CODEC
output reg LRCLK;			// Left/Right clock to CODEC
output reg SDin;			// forms serial data in to CODEC
input SDout;			// from CODEC SDout pin (serial data in to core)
output reg AMP_ON;			// signal to turn amp on
output reg RSTn;			// active low reset to CODEC

wire rst_n;				// internal global active low reset
wire valid;
wire strt_cnv,cnv_cmplt,valid_fall,valid_rise;
wire [15:0] lft_in,rht_in;
wire [15:0] lft_out,rht_out,lft_out_sel,rht_out_sel;
wire [2:0] chnnl;
wire [11:0] res;
wire [11:0] LP_gain,B1_gain,B2_gain,B3_gain,HP_gain,volume;


reg [10:0] del;

/////////////////////////////////////
// Instantiate Reset synchronizer //
///////////////////////////////////
//rst_synch iRST(.clk(clk),.RST_n(RST_n),.rst_n(rst_n));

			  
///////////////////////////////////////////
// Instantiate Your Slide Pot Interface //
/////////////////////////////////////////
slide_intf iSLD(.POT_LP(LP_gain), .POT_B1(B1_gain), .POT_B2(B2_gain), .POT_B3(B3_gain), 
                .POT_HP(HP_gain), .VOLUME(volume),.MISO(A2D_MISO),.MOSI(A2D_MOSI),
             .SCLK(A2D_SCLK),.clk(clk),.rst_n(RST_n),.a2d_SS_n(A2D_SS_n));
	
				
///////////////////////////////////////
// Instantiate Your CODEC Interface //
/////////////////////////////////////
//codec_intf iCS(.clk(clk), .rst_n(rst_n), .lft_in(lft_in), .rht_in(rht_in), .lft_out(lft_out), .rht_out(rht_out),
//                  .valid(valid), .RSTn(RSTn), .MCLK(MCLK), .SCLK(SCL), .LRCLK(LRCLK), .SDin(SDin), .SDout(SDout));
//
///////////////////////////////////
// Instantiate Equalizer Engine //
/////////////////////////////////
dig_core_intf iDig(.clk(clk), .rst_n(rst_n), .lft_in(lft_in), .rht_in(rht_in), .lft_out(lft_out), .rht_out(rht_out), 
		.valid(valid), .POT_B1(B1_gain),.POT_B2(B2_gain), .POT_B3(B3_gain), .POT_HP(HP_gain), .POT_LP(LP_gain),
		 .POT_VOL(volume), .AMP_ON(AMP_ON));
EqualizerLoopBack iLoop(.clk(clk), .RST_n(RST_n), .SDin(SDin), .SDout(SDout), .RSTn(RSTn), .SCL(SCL), .MCLK(MCLK), .LRCLK(LRCLK));


////////////////////////////////////////////////////////////
// Instantiate LED effect driver (optional extra credit) //
//////////////////////////////////////////////////////////
assign LED  = (volume < 64) ? 8'h00 :
	      (volume <=1024) ? 8'h01:
	      (volume <= 2048) ? 8'h03:
	      (volume <= 3072) ? 8'h07:
	      (volume <= 4096) ? 8'h0f:
	      (volume <= 5120) ? 8'h1f:
	      (volume <= 6144) ? 8'h3f:
	      (volume <= 7168) ? 8'h7f: 8'hff;
///////////////////////////////////////////////
// Implement logic for delaying Amp on till //
// after queues are steady.   (AMP_ON)     //
////////////////////////////////////////////
//done in dig_core_intf


endmodule
